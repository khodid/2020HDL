module module RANDOM_CNT (nRST, CLK, CLR, EN, UP_DOWN, JUMP_NUM, CNTo);

endmodule // module RANDOM_CNT (nRST, CLK, CLR, EN, UP_DOWN, JUMP_NUM, CNTo);
