module module DATA_ORDER(nRST, CLK, DATAi, VALi, MAX1st, MAX2nd, MAX3rd, MIN1st,
MIN2nd, MIN3rd, AVEo);

endmodule // module DATA_ORDER(nRST, CLK, DATAi, VALi, MAX1st, MAX2nd, MAX3rd, MIN1st,
MIN2nd, MIN3rd, AVEo);
